module testbench();

	timeunit 10ns;
	timeprecision 1ns;
	
	logic [7:0] A,B,S;
	logic X;
	logic [16:0] Sol;
	
	



endmodule 