/*module multiply ( 
	input logic [7:0] B, S,
	input logic X, 
	output logic [7:0] A,
	
);

always_comb begin	
	case (B[0])
		1'b0 : begin
			shift bitshift (asdfasdf);
		end
		1'b1 : begin
			ripple_adder asdf (.A(), .B(), .cin(), .S(), .cout());
			shift bitshift1 (asdfasdf);
		end
	endcase
end
















endmodules
*/